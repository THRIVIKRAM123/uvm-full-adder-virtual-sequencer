class v_seqr extends uvm_sequencer#(xtn);
	`uvm_component_utils(v_seqr)
	
              seqr seqr_h;

          function new(string name = "v_seqr", uvm_component parent = null);
    super.new(name, parent);
  endfunction

	

endclass